library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 10
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture rtl of rom is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);
  
  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
        -- Inicializa os endereços:
--        tmp(0) := "0000" & "000" & "000000000"; -- Load for r7 mem [0x200]
--        tmp(1) := "0000" & "000" & "000000000"; -- Jump to line of the code [256]
--        tmp(2) := "0000" & "000" & "000000000";
--        tmp(3) := "0110" & "000" & "000000110"; -- JUMP
--        tmp(4) := "0000" & "000" & "000000000";
--        tmp(5) := "0000" & "000" & "000000000";
--        tmp(6) := "0000" & "000" & "000000000";
--        tmp(7) := "0111" & "000" & "000000010"; -- JE
--        tmp(8) := "0000" & "000" & "000000000";
--        tmp(9) := "0000" & "000" & "000000000";
--        tmp(10) := "0000" & "000" & "000000000";
--        tmp(256) := x"55";
--        tmp(0) := "0000" & "000" & "000000000"; -- 
--        tmp(1) := "0000" & "000" & "000000000"; -- 
		  -- CMP
--        tmp(2) := "0001" & "001" & "000001111"; -- LOAD R1, #15
--        tmp(3) := "0000" & "000" & "000000000"; -- NOP
--        tmp(4) := "1000" & "001" & "010000011"; -- STORE Mem[131], R1
--        tmp(5) := "1001" & "001" & "010000011"; -- CMP R1, Mem[131]
--        tmp(6) := "0111" & "000" & "000001001"; -- JE ROM[9]
			-- ADD
--        tmp(2) := "0001" & "001" & "000001111"; -- LOAD R1, #15
--		  tmp(3) := "0001" & "010" & "000011110"; -- LOAD R1, #30
--        tmp(4) := "0000" & "000" & "000000000"; -- NOP
--        tmp(5) := "1000" & "001" & "010000011"; -- STORE Mem[131], R1
--		  tmp(6) := "1000" & "010" & "010000111"; -- STORE Mem[131], R1
--        tmp(7) := "0010" & "001" & "010000011"; -- ADD R1, Mem[131]
--        tmp(8) := "1001" & "001" & "010000111"; -- CMP R1, Mem[135]
--        tmp(9) := "0111" & "000" & "000000000"; -- JE ROM[0]
--        tmp(10) := "0000" & "000" & "000000000"; -- NOP
--        tmp(11) := "0000" & "000" & "000000000"; -- NOP
--        tmp(12) := "0110" & "000" & "000000000"; -- JUMP
--		  -- SUB
--        tmp(2) := "0001" & "001" & "000001111"; -- LOAD R1, #15
--		  tmp(3) := "0001" & "010" & "000000000"; -- LOAD R1, #0
--        tmp(4) := "0000" & "000" & "000000000"; -- NOP
--        tmp(5) := "1000" & "001" & "010000011"; -- STORE Mem[131], R1
--		  tmp(6) := "1000" & "010" & "010000111"; -- STORE Mem[135], R1
--        tmp(7) := "0011" & "001" & "010000011"; -- SUB R1, Mem[131]
--        tmp(8) := "1001" & "001" & "010000111"; -- CMP R1, Mem[135]
--        tmp(9) := "0111" & "000" & "000000000"; -- JE ROM[9]
--        tmp(10) := "0000" & "000" & "000000000"; -- JE ROM[9]
--        tmp(11) := "0000" & "000" & "000000000"; -- JE ROM[9]
--        tmp(12) := "0110" & "000" & "000000000"; -- JUMP
-- STORE ON IO
--        tmp(2) := "0001" & "001" & "000000010"; -- LOAD R1, #2
--		  tmp(3) := "0001" & "010" & "000000001"; -- LOAD R2, #1
--        tmp(4) := "0000" & "000" & "000000000"; -- NOP
--        tmp(5) := "1000" & "001" & "010000011"; -- STORE Mem[131], R1
--		  tmp(6) := "1000" & "010" & "010000111"; -- STORE Mem[135], R1
--        tmp(7) := "0010" & "001" & "010000011"; -- ADD R1, Mem[131]
--		  tmp(8) := "1000" & "001" & "000000000"; -- STORE R1, Mem[0]
--        tmp(9) := "0110" & "000" & "000000111"; -- JUMP

-- ADDI
--        tmp(2) := "0001" & "001" & "000001111"; -- LOAD R1, #15
--		  tmp(3) := "0001" & "010" & "000010000"; -- LOAD R2, #16
--        tmp(4) := "0000" & "000" & "000000000"; -- NOP
--        tmp(5) := "1000" & "001" & "010000011"; -- STORE Mem[131], R1
--		  tmp(6) := "1000" & "010" & "010000111"; -- STORE Mem[135], R2
--        tmp(7) := "0010" & "001" & "000000001"; -- ADDI R1, #1
--        tmp(8) := "1001" & "001" & "010000111"; -- CMP R1, Mem[135]
--        tmp(9) := "0111" & "000" & "000000000"; -- JE ROM[9]
--        tmp(10) := "0000" & "000" & "000000000"; -- NOP
--        tmp(11) := "0000" & "000" & "000000000"; -- NOP
--        tmp(12) := "0110" & "000" & "000000000"; -- JUMP

-- TESTE ZERANDO R1

--tmp(0) := "0001000000000000"; -- LOAD R0, #0
--tmp(1) := "1000000000000000"; -- STORE R0, %0
--tmp(2) := "0001001000000001"; -- LOAD R1, #1
--tmp(3) := "1000001000000001"; -- STORE R1, %1
--tmp(4) := "0001010000000010"; -- LOAD R2, #2
--tmp(5) := "1000010000000010"; -- STORE R2, %2
--tmp(6) := "0001000000000011"; -- LOAD R0, #3
--tmp(7) := "0010000000000001"; -- ADD R0, %1
--tmp(8) := "1000000000000011"; -- STORE R0, %3
--tmp(9) := "0001000000000000"; -- LOAD R0, #0
--tmp(10) := "0010000000001111"; -- ADD R0, %15
--tmp(11) := "1000000000000100"; -- STORE R0, %4
--tmp(12) := "0001000000000000"; -- LOAD R0, #0
--tmp(13) := "0010000000010000"; -- ADD R0, %16
--tmp(14) := "1000000000000101"; -- STORE R0, %5

--tmp(0) := "0001000000000000"; -- LOAD R0, #0
--tmp(1) := "1000000000000000"; -- STORE R0, %0
--tmp(2) := "1000000000000001"; -- STORE R0, %1
--tmp(3) := "1000000000000010"; -- STORE R0, %2
--tmp(4) := "1000000000000011"; -- STORE R0, %3
--tmp(5) := "1000000000000100"; -- STORE R0, %4
--tmp(6) := "1000000000000101"; -- STORE R0, %5
--tmp(7) := "0001000000000000"; -- LOOP: LOAD R0, #0
--tmp(8) := "1001000000001111"; -- CMP R0, %15
--tmp(9) := "0111000000000111"; -- JE LOOP
--tmp(10) := "0001001000000000"; -- LOAD R1, #0
--tmp(11) := "1000001000010000"; -- STORE R1, %16
--tmp(12) := "0001001000000001"; -- LOAD R1, #1
--tmp(13) := "0010001000000000"; -- ADD R1, %0
--tmp(14) := "1000001000000000"; -- STORE R1, %0
--tmp(15) := "0001010000001010"; -- IFS: LOAD R2, #10
--tmp(16) := "1001010000000000"; -- CMP R2, %0
--tmp(17) := "0111000000100010"; -- JE INC_SEC_D
--tmp(18) := "0001010000000110"; -- LOAD R2, #6
--tmp(19) := "1001010000000001"; -- CMP R2, %1
--tmp(20) := "0111000000101000"; -- JE INC_MIN_U
--tmp(21) := "0001010000001010"; -- LOAD R2, #10
--tmp(22) := "1001010000000010"; -- CMP R2, %2
--tmp(23) := "0111000000101110"; -- JE INC_MIN_D
--tmp(24) := "0001010000000110"; -- LOAD R2, #6
--tmp(25) := "1001010000000011"; -- CMP R2, %3
--tmp(26) := "0111000000110100"; -- JE INC_HOUR_U
--tmp(27) := "0001010000001010"; -- LOAD R2, #10
--tmp(28) := "1001010000000100"; -- CMP R2, %4
--tmp(29) := "0111000000111010"; -- JE INC_HOUR_D
--tmp(30) := "0001010000000010"; -- LOAD R2, #2
--tmp(31) := "1001010000000101"; -- CMP R2, %5
--tmp(32) := "0111000001000000"; -- JE DAY
--tmp(33) := "0110000000000111"; -- JMP LOOP
--tmp(34) := "0001001000000001"; -- INC_SEC_D: LOAD R1, #1
--tmp(35) := "0010001000000001"; -- ADD R1, %1
--tmp(36) := "1000001000000001"; -- STORE R1, %1
--tmp(37) := "0001000000000000"; -- LOAD R0, #0
--tmp(38) := "1000000000000000"; -- STORE R0, %0
--tmp(39) := "0110000000001111"; -- JMP IFS
--tmp(40) := "0001001000000001"; -- INC_MIN_U: LOAD R1, #1
--tmp(41) := "0010001000000010"; -- ADD R1, %2
--tmp(42) := "1000001000000010"; -- STORE R1, %2
--tmp(43) := "0001000000000000"; -- LOAD R0, #0
--tmp(44) := "1000000000000001"; -- STORE R0, %1
--tmp(45) := "0110000000001111"; -- JMP IFS
--tmp(46) := "0001001000000001"; -- INC_MIN_D: LOAD R1, #1
--tmp(47) := "0010001000000011"; -- ADD R1, %3
--tmp(48) := "1000001000000011"; -- STORE R1, %3
--tmp(49) := "0001000000000000"; -- LOAD R0, #0
--tmp(50) := "1000000000000010"; -- STORE R0, %2
--tmp(51) := "0110000000001111"; -- JMP IFS
--tmp(52) := "0001001000000001"; -- INC_HOUR_U: LOAD R1, #1
--tmp(53) := "0010001000000100"; -- ADD R1, %4
--tmp(54) := "1000001000000100"; -- STORE R1, %4
--tmp(55) := "0001000000000000"; -- LOAD R0, #0
--tmp(56) := "1000000000000011"; -- STORE R0, %3
--tmp(57) := "0110000000001111"; -- JMP IFS
--tmp(58) := "0001001000000001"; -- INC_HOUR_D: LOAD R1, #1
--tmp(59) := "0010001000000101"; -- ADD R1, %5
--tmp(60) := "1000001000000101"; -- STORE R1, %5
--tmp(61) := "0001000000000000"; -- LOAD R0, #0
--tmp(62) := "1000000000000100"; -- STORE R0, %4
--tmp(63) := "0110000000001111"; -- JMP IFS
--tmp(64) := "0001001000000100"; -- DAY: LOAD R1, #4
--tmp(65) := "1001001000000100"; -- CMP R1, %4
--tmp(66) := "0111000001000100"; -- JE RESET_DAY
--tmp(67) := "0110000000000111"; -- JMP LOOP
--tmp(68) := "0001000000000000"; -- RESET_DAY: LOAD R0, #0
--tmp(69) := "1000000000000000"; -- STORE R0, %0
--tmp(70) := "1000000000000001"; -- STORE R0, %1
--tmp(71) := "1000000000000010"; -- STORE R0, %2
--tmp(72) := "1000000000000011"; -- STORE R0, %3
--tmp(73) := "1000000000000100"; -- STORE R0, %4
--tmp(74) := "1000000000000101"; -- STORE R0, %5
--tmp(75) := "0110000000000111"; -- JMP LOOP

--tmp(0) := "0001000000000000"; -- LOAD R0, #0
--tmp(1) := "1000000000000000"; -- STORE R0, %0
--tmp(2) := "1000000000000001"; -- STORE R0, %1
--tmp(3) := "1000000000000010"; -- STORE R0, %2
--tmp(4) := "1000000000000011"; -- STORE R0, %3
--tmp(5) := "1000000000000100"; -- STORE R0, %4
--tmp(6) := "1000000000000101"; -- STORE R0, %5
--tmp(7) := "1000000010000010"; -- STORE R0, %130
--tmp(8) := "1000000010000011"; -- STORE R0, %131
--tmp(9) := "1000000010000100"; -- STORE R0, %132
--tmp(10) := "1000000010000101"; -- STORE R0, %133
--tmp(11) := "1000000010000110"; -- STORE R0, %134
--tmp(12) := "1000000010000111"; -- STORE R0, %135
--tmp(13) := "0001001000000001"; -- LOAD R1, #1
--tmp(14) := "1000001000010000"; -- STORE R1, %16
--tmp(15) := "0001000000000000"; -- LOOP: LOAD R0, #0
--tmp(16) := "1001000000001111"; -- CMP R0, %15
--tmp(17) := "0111000000001111"; -- JE LOOP
--tmp(18) := "0001001000000001"; -- LOAD R1, #1
--tmp(19) := "1000001000010000"; -- STORE R1, %16
--tmp(20) := "0001001000000001"; -- LOAD R1, #1
--tmp(21) := "0010001010000010"; -- ADD R1, %130
--tmp(22) := "1000001000000000"; -- STORE R1, %0
--tmp(23) := "1000001010000010"; -- STORE R1, %130
--tmp(24) := "0001010000001010"; -- IFS: LOAD R2, #10
--tmp(25) := "1001010010000010"; -- CMP R2, %130
--tmp(26) := "0111000000101011"; -- JE INC_SEC_D
--tmp(27) := "0001010000000110"; -- LOAD R2, #6
--tmp(28) := "1001010010000011"; -- CMP R2, %131
--tmp(29) := "0111000000110011"; -- JE INC_MIN_U
--tmp(30) := "0001010000001010"; -- LOAD R2, #10
--tmp(31) := "1001010010000100"; -- CMP R2, %132
--tmp(32) := "0111000000111011"; -- JE INC_MIN_D
--tmp(33) := "0001010000000110"; -- LOAD R2, #6
--tmp(34) := "1001010010000101"; -- CMP R2, %133
--tmp(35) := "0111000001000011"; -- JE INC_HOUR_U
--tmp(36) := "0001010000001010"; -- LOAD R2, #10
--tmp(37) := "1001010010000110"; -- CMP R2, %134
--tmp(38) := "0111000001001011"; -- JE INC_HOUR_D
--tmp(39) := "0001010000000010"; -- LOAD R2, #2
--tmp(40) := "1001010010000111"; -- CMP R2, %135
--tmp(41) := "0111000001010011"; -- JE DAY
--tmp(42) := "0110000000001111"; -- JMP LOOP
--tmp(43) := "0001001000000001"; -- INC_SEC_D: LOAD R1, #1
--tmp(44) := "0010001010000011"; -- ADD R1, %131
--tmp(45) := "1000001010000011"; -- STORE R1, %131
--tmp(46) := "1000001000000001"; -- STORE R1, %1
--tmp(47) := "0001000000000000"; -- LOAD R0, #0
--tmp(48) := "1000000010000010"; -- STORE R0, %130
--tmp(49) := "1000000000000000"; -- STORE R0, %0
--tmp(50) := "0110000000011000"; -- JMP IFS
--tmp(51) := "0001001000000001"; -- INC_MIN_U: LOAD R1, #1
--tmp(52) := "0010001010000100"; -- ADD R1, %132
--tmp(53) := "1000001010000100"; -- STORE R1, %132
--tmp(54) := "1000001000000010"; -- STORE R1, %2
--tmp(55) := "0001000000000000"; -- LOAD R0, #0
--tmp(56) := "1000000010000011"; -- STORE R0, %131
--tmp(57) := "1000000000000001"; -- STORE R0, %1
--tmp(58) := "0110000000011000"; -- JMP IFS
--tmp(59) := "0001001000000001"; -- INC_MIN_D: LOAD R1, #1
--tmp(60) := "0010001010000101"; -- ADD R1, %133
--tmp(61) := "1000001010000101"; -- STORE R1, %133
--tmp(62) := "1000001000000011"; -- STORE R1, %3
--tmp(63) := "0001000000000000"; -- LOAD R0, #0
--tmp(64) := "1000000010000100"; -- STORE R0, %132
--tmp(65) := "1000000000000010"; -- STORE R0, %2
--tmp(66) := "0110000000011000"; -- JMP IFS
--tmp(67) := "0001001000000001"; -- INC_HOUR_U: LOAD R1, #1
--tmp(68) := "0010001010000110"; -- ADD R1, %134
--tmp(69) := "1000001010000110"; -- STORE R1, %134
--tmp(70) := "1000001000000100"; -- STORE R1, %4
--tmp(71) := "0001000000000000"; -- LOAD R0, #0
--tmp(72) := "1000000010000101"; -- STORE R0, %133
--tmp(73) := "1000000000000011"; -- STORE R0, %3
--tmp(74) := "0110000000011000"; -- JMP IFS
--tmp(75) := "0001001000000001"; -- INC_HOUR_D: LOAD R1, #1
--tmp(76) := "0010001010000111"; -- ADD R1, %135
--tmp(77) := "1000001010000111"; -- STORE R1, %135
--tmp(78) := "1000001000000101"; -- STORE R1, %5
--tmp(79) := "0001000000000000"; -- LOAD R0, #0
--tmp(80) := "1000000010000110"; -- STORE R0, %134
--tmp(81) := "1000000000000100"; -- STORE R0, %4
--tmp(82) := "0110000000011000"; -- JMP IFS
--tmp(83) := "0001001000000100"; -- DAY: LOAD R1, #4
--tmp(84) := "1001001010000110"; -- CMP R1, %134
--tmp(85) := "0111000001010111"; -- JE RESET_DAY
--tmp(86) := "0110000000001111"; -- JMP LOOP
--tmp(87) := "0001000000000000"; -- RESET_DAY: LOAD R0, #0
--tmp(88) := "1000000000000000"; -- STORE R0, %0
--tmp(89) := "1000000000000001"; -- STORE R0, %1
--tmp(90) := "1000000000000010"; -- STORE R0, %2
--tmp(91) := "1000000000000011"; -- STORE R0, %3
--tmp(92) := "1000000000000100"; -- STORE R0, %4
--tmp(93) := "1000000000000101"; -- STORE R0, %5
--tmp(94) := "1000000010000010"; -- STORE R0, %130
--tmp(95) := "1000000010000011"; -- STORE R0, %131
--tmp(96) := "1000000010000100"; -- STORE R0, %132
--tmp(97) := "1000000010000101"; -- STORE R0, %133
--tmp(98) := "1000000010000110"; -- STORE R0, %134
--tmp(99) := "1000000010000111"; -- STORE R0, %135
--tmp(100) := "0110000000001111"; -- JMP LOOP

	tmp(0) := "0001000000000000"; -- LOAD R0, #0
	tmp(1) := "1000000000000000"; -- STORE R0, %0
	tmp(2) := "1000000000000001"; -- STORE R0, %1
	tmp(3) := "1000000000000010"; -- STORE R0, %2
	tmp(4) := "1000000000000011"; -- STORE R0, %3
	tmp(5) := "1000000000000100"; -- STORE R0, %4
	tmp(6) := "1000000000000101"; -- STORE R0, %5
	tmp(7) := "1000000010000010"; -- STORE R0, %130
	tmp(8) := "1000000010000011"; -- STORE R0, %131
	tmp(9) := "1000000010000100"; -- STORE R0, %132
	tmp(10) := "1000000010000101"; -- STORE R0, %133
	tmp(11) := "1000000010000110"; -- STORE R0, %134
	tmp(12) := "1000000010000111"; -- STORE R0, %135
	tmp(13) := "0001001000000001"; -- LOAD R1, #1
	tmp(14) := "1000001000010000"; -- STORE R1, %16
	tmp(15) := "0001000000000000"; -- LOOP: LOAD R0, #0
	tmp(16) := "1001000000001111"; -- CMP R0, %15
	tmp(17) := "0111000000001111"; -- JE LOOP
	tmp(18) := "0001001000000001"; -- LOAD R1, #1
	tmp(19) := "1000001000010000"; -- STORE R1, %16
	tmp(20) := "0001010000000010"; -- LOAD R2, #2
	tmp(21) := "1001010000000110"; -- CMP R2, %6
	tmp(22) := "0111000001101110"; -- JE CONFIG_SEC
	tmp(23) := "0001010000000100"; -- LOAD R2, #4
	tmp(24) := "1001010000000110"; -- CMP R2, %6
	tmp(25) := "0111000010000101"; -- JE CONFIG_MIN
	tmp(26) := "0001010000001000"; -- LOAD R2, #8
	tmp(27) := "1001010000000110"; -- CMP R2, %6
	tmp(28) := "0111000010011100"; -- JE CONFIG_HOUR
	tmp(29) := "0001001000000001"; -- LOAD R1, #1
	tmp(30) := "0010001010000010"; -- ADD R1, %130
	tmp(31) := "1000001000000000"; -- STORE R1, %0
	tmp(32) := "1000001010000010"; -- STORE R1, %130
	tmp(33) := "0001010000001010"; -- IFS: LOAD R2, #10
	tmp(34) := "1001010010000010"; -- CMP R2, %130
	tmp(35) := "0111000000110100"; -- JE INC_SEC_D
	tmp(36) := "0001010000000110"; -- LOAD R2, #6
	tmp(37) := "1001010010000011"; -- CMP R2, %131
	tmp(38) := "0111000000111100"; -- JE INC_MIN_U
	tmp(39) := "0001010000001010"; -- LOAD R2, #10
	tmp(40) := "1001010010000100"; -- CMP R2, %132
	tmp(41) := "0111000001000100"; -- JE INC_MIN_D
	tmp(42) := "0001010000000110"; -- LOAD R2, #6
	tmp(43) := "1001010010000101"; -- CMP R2, %133
	tmp(44) := "0111000001001100"; -- JE INC_HOUR_U
	tmp(45) := "0001010000001010"; -- LOAD R2, #10
	tmp(46) := "1001010010000110"; -- CMP R2, %134
	tmp(47) := "0111000001010100"; -- JE INC_HOUR_D
	tmp(48) := "0001010000000010"; -- LOAD R2, #2
	tmp(49) := "1001010010000111"; -- CMP R2, %135
	tmp(50) := "0111000001011100"; -- JE DAY
	tmp(51) := "0110000000001111"; -- JMP LOOP
	tmp(52) := "0001001000000001"; -- INC_SEC_D: LOAD R1, #1
	tmp(53) := "0010001010000011"; -- ADD R1, %131
	tmp(54) := "1000001010000011"; -- STORE R1, %131
	tmp(55) := "1000001000000001"; -- STORE R1, %1
	tmp(56) := "0001000000000000"; -- LOAD R0, #0
	tmp(57) := "1000000010000010"; -- STORE R0, %130
	tmp(58) := "1000000000000000"; -- STORE R0, %0
	tmp(59) := "0110000000100001"; -- JMP IFS
	tmp(60) := "0001001000000001"; -- INC_MIN_U: LOAD R1, #1
	tmp(61) := "0010001010000100"; -- ADD R1, %132
	tmp(62) := "1000001010000100"; -- STORE R1, %132
	tmp(63) := "1000001000000010"; -- STORE R1, %2
	tmp(64) := "0001000000000000"; -- LOAD R0, #0
	tmp(65) := "1000000010000011"; -- STORE R0, %131
	tmp(66) := "1000000000000001"; -- STORE R0, %1
	tmp(67) := "0110000000100001"; -- JMP IFS
	tmp(68) := "0001001000000001"; -- INC_MIN_D: LOAD R1, #1
	tmp(69) := "0010001010000101"; -- ADD R1, %133
	tmp(70) := "1000001010000101"; -- STORE R1, %133
	tmp(71) := "1000001000000011"; -- STORE R1, %3
	tmp(72) := "0001000000000000"; -- LOAD R0, #0
	tmp(73) := "1000000010000100"; -- STORE R0, %132
	tmp(74) := "1000000000000010"; -- STORE R0, %2
	tmp(75) := "0110000000100001"; -- JMP IFS
	tmp(76) := "0001001000000001"; -- INC_HOUR_U: LOAD R1, #1
	tmp(77) := "0010001010000110"; -- ADD R1, %134
	tmp(78) := "1000001010000110"; -- STORE R1, %134
	tmp(79) := "1000001000000100"; -- STORE R1, %4
	tmp(80) := "0001000000000000"; -- LOAD R0, #0
	tmp(81) := "1000000010000101"; -- STORE R0, %133
	tmp(82) := "1000000000000011"; -- STORE R0, %3
	tmp(83) := "0110000000100001"; -- JMP IFS
	tmp(84) := "0001001000000001"; -- INC_HOUR_D: LOAD R1, #1
	tmp(85) := "0010001010000111"; -- ADD R1, %135
	tmp(86) := "1000001010000111"; -- STORE R1, %135
	tmp(87) := "1000001000000101"; -- STORE R1, %5
	tmp(88) := "0001000000000000"; -- LOAD R0, #0
	tmp(89) := "1000000010000110"; -- STORE R0, %134
	tmp(90) := "1000000000000100"; -- STORE R0, %4
	tmp(91) := "0110000000100001"; -- JMP IFS
	tmp(92) := "0001001000000100"; -- DAY: LOAD R1, #4
	tmp(93) := "1001001010000110"; -- CMP R1, %134
	tmp(94) := "0111000001100000"; -- JE RESET_DAY
	tmp(95) := "0110000000001111"; -- JMP LOOP
	tmp(96) := "0001000000000000"; -- RESET_DAY: LOAD R0, #0
	tmp(97) := "1000000000000000"; -- STORE R0, %0
	tmp(98) := "1000000000000001"; -- STORE R0, %1
	tmp(99) := "1000000000000010"; -- STORE R0, %2
	tmp(100) := "1000000000000011"; -- STORE R0, %3
	tmp(101) := "1000000000000100"; -- STORE R0, %4
	tmp(102) := "1000000000000101"; -- STORE R0, %5
	tmp(103) := "1000000010000010"; -- STORE R0, %130
	tmp(104) := "1000000010000011"; -- STORE R0, %131
	tmp(105) := "1000000010000100"; -- STORE R0, %132
	tmp(106) := "1000000010000101"; -- STORE R0, %133
	tmp(107) := "1000000010000110"; -- STORE R0, %134
	tmp(108) := "1000000010000111"; -- STORE R0, %135
	tmp(109) := "0110000000001111"; -- JMP LOOP
	tmp(110) := "0001001000000001"; -- CONFIG_SEC: LOAD R1, #1
	tmp(111) := "0010001010000010"; -- ADD R1, %130
	tmp(112) := "1000001000000000"; -- STORE R1, %0
	tmp(113) := "1000001010000010"; -- STORE R1, %130
	tmp(114) := "0001010000001010"; -- CONFIG_SEC_IF: LOAD R2, #10
	tmp(115) := "1001010010000010"; -- CMP R2, %130
	tmp(116) := "0111000001111001"; -- JE CONFIG_INC_SEC_D
	tmp(117) := "0001010000000110"; -- LOAD R2, #6
	tmp(118) := "1001010010000011"; -- CMP R2, %131
	tmp(119) := "0111000010000001"; -- JE CONFIG_RESET_SEC_D
	tmp(120) := "0110000000001111"; -- JMP LOOP
	tmp(121) := "0001001000000001"; -- CONFIG_INC_SEC_D: LOAD R1, #1
	tmp(122) := "0010001010000011"; -- ADD R1, %131
	tmp(123) := "1000001010000011"; -- STORE R1, %131
	tmp(124) := "1000001000000001"; -- STORE R1, %1
	tmp(125) := "0001000000000000"; -- LOAD R0, #0
	tmp(126) := "1000000010000010"; -- STORE R0, %130
	tmp(127) := "1000000000000000"; -- STORE R0, %0
	tmp(128) := "0110000001110010"; -- JMP CONFIG_SEC_IF
	tmp(129) := "0001000000000000"; -- CONFIG_RESET_SEC_D: LOAD R0, #0
	tmp(130) := "1000000010000011"; -- STORE R0, %131
	tmp(131) := "1000000000000001"; -- STORE R0, %1
	tmp(132) := "0110000000001111"; -- JMP LOOP
	tmp(133) := "0001001000000001"; -- CONFIG_MIN: LOAD R1, #1
	tmp(134) := "0010001010000100"; -- ADD R1, %132
	tmp(135) := "1000001010000100"; -- STORE R1, %132
	tmp(136) := "1000001000000010"; -- STORE R1, %2
	tmp(137) := "0001010000001010"; -- CONFIG_MIN_IF: LOAD R2, #10
	tmp(138) := "1001010010000100"; -- CMP R2, %132
	tmp(139) := "0111000010010000"; -- JE CONFIG_INC_MIN_D
	tmp(140) := "0001010000000110"; -- LOAD R2, #6
	tmp(141) := "1001010010000101"; -- CMP R2, %133
	tmp(142) := "0111000010011000"; -- JE CONFIG_RESET_MIN_D
	tmp(143) := "0110000000001111"; -- JMP LOOP
	tmp(144) := "0001001000000001"; -- CONFIG_INC_MIN_D: LOAD R1, #1
	tmp(145) := "0010001010000101"; -- ADD R1, %133
	tmp(146) := "1000001010000101"; -- STORE R1, %133
	tmp(147) := "1000001000000011"; -- STORE R1, %3
	tmp(148) := "0001000000000000"; -- LOAD R0, #0
	tmp(149) := "1000000010000100"; -- STORE R0, %132
	tmp(150) := "1000000000000010"; -- STORE R0, %2
	tmp(151) := "0110000010001001"; -- JMP CONFIG_MIN_IF
	tmp(152) := "0001000000000000"; -- CONFIG_RESET_MIN_D: LOAD R0, #0
	tmp(153) := "1000000010000101"; -- STORE R0, %133
	tmp(154) := "1000000000000011"; -- STORE R0, %3
	tmp(155) := "0110000000001111"; -- JMP LOOP
	tmp(156) := "0001001000000001"; -- CONFIG_HOUR: LOAD R1, #1
	tmp(157) := "0010001010000110"; -- ADD R1, %134
	tmp(158) := "1000001010000110"; -- STORE R1, %134
	tmp(159) := "1000001000000100"; -- STORE R1, %4
	tmp(160) := "0001010000001010"; -- CONFIG_HOUR_IF: LOAD R2, #10
	tmp(161) := "1001010010000110"; -- CMP R2, %134
	tmp(162) := "0111000010100111"; -- JE CONFIG_INC_HOUR_D
	tmp(163) := "0001010000000010"; -- LOAD R2, #2
	tmp(164) := "1001010010000111"; -- CMP R2, %135
	tmp(165) := "0111000010101111"; -- JE CONFIG_DAY
	tmp(166) := "0110000000001111"; -- JMP LOOP
	tmp(167) := "0001001000000001"; -- CONFIG_INC_HOUR_D: LOAD R1, #1
	tmp(168) := "0010001010000111"; -- ADD R1, %135
	tmp(169) := "1000001010000111"; -- STORE R1, %135
	tmp(170) := "1000001000000101"; -- STORE R1, %5
	tmp(171) := "0001000000000000"; -- LOAD R0, #0
	tmp(172) := "1000000010000110"; -- STORE R0, %134
	tmp(173) := "1000000000000100"; -- STORE R0, %4
	tmp(174) := "0110000010100000"; -- JMP CONFIG_HOUR_IF
	tmp(175) := "0001001000000100"; -- CONFIG_DAY: LOAD R1, #4
	tmp(176) := "1001001010000110"; -- CMP R1, %134
	tmp(177) := "0111000010110011"; -- JE CONFIG_RESET_DAY
	tmp(178) := "0110000000001111"; -- JMP LOOP
	tmp(179) := "0001000000000000"; -- CONFIG_RESET_DAY: LOAD R0, #0
	tmp(180) := "1000000000000100"; -- STORE R0, %4
	tmp(181) := "1000000000000101"; -- STORE R0, %5
	tmp(182) := "1000000010000110"; -- STORE R0, %134
	tmp(183) := "1000000010000111"; -- STORE R0, %135
	tmp(184) := "0110000000001111"; -- JMP LOOP
       return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;